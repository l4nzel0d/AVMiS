library verilog;
use verilog.vl_types.all;
entity pract1_vlg_vec_tst is
end pract1_vlg_vec_tst;
