library verilog;
use verilog.vl_types.all;
entity pract5_vlg_vec_tst is
end pract5_vlg_vec_tst;
