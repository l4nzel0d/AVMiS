library verilog;
use verilog.vl_types.all;
entity pract4 is
    port(
        X2              : in     vl_logic;
        X1              : in     vl_logic;
        X0              : in     vl_logic;
        E               : in     vl_logic;
        Y0              : out    vl_logic;
        Y1              : out    vl_logic;
        Y2              : out    vl_logic;
        Y3              : out    vl_logic;
        Y4              : out    vl_logic;
        Y5              : out    vl_logic;
        Y6              : out    vl_logic;
        Y7              : out    vl_logic
    );
end pract4;
