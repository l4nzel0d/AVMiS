library verilog;
use verilog.vl_types.all;
entity pract4_vlg_vec_tst is
end pract4_vlg_vec_tst;
