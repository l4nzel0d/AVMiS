library verilog;
use verilog.vl_types.all;
entity pract6_vlg_vec_tst is
end pract6_vlg_vec_tst;
